module submodule(
    input a,
    output b
);

assign b = ~a;

endmodule